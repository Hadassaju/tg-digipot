magic
tech sky130A
timestamp 1698428228
<< end >>
