** sch_path: /foss/designs/tg-tb.sch
**.subckt tg-tb
Vdd vd GND 1.8
.save i(vdd)
Vin in GND pulse 0 1.8 '0.495/ 1 ' '0.01/1 ' '0.01/1 ' '0.49/1 ' '1/1 '
x1 vd in GND A B tg
Va A GND 0.9
.save i(va)
C1 net1 net2 1p m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.control
save all
tran 1m 3
let Vab = V(A)-V(B)
let R = Vab/i(Va)
plot abs(R)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/tg.sym # of pins=5
** sym_path: /foss/designs/tg.sym
** sch_path: /foss/designs/tg.sch
.subckt tg vd ctrl vgnd A B
*.iopin B
*.iopin A
*.iopin vgnd
*.iopin vd
*.ipin ctrl
x1 vd ctrl nctrl vgnd inverter
XM1 A ctrl B vgnd sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 A nctrl B vd sky130_fd_pr__pfet_01v8 L=0.15 W=30 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/inverter/xschem_files/inverter.sym # of pins=4
** sym_path: /foss/designs/inverter/xschem_files/inverter.sym
** sch_path: /foss/designs/inverter/xschem_files/inverter.sch
.subckt inverter vd in out gnd
*.ipin in
*.opin out
*.iopin vd
*.iopin gnd
XN0 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XP0 out in vd vd sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
