magic
tech sky130A
magscale 1 2
timestamp 1698427088
<< error_p >>
rect 19 231 77 237
rect 19 197 31 231
rect 19 191 77 197
rect -77 -197 -19 -191
rect -77 -231 -65 -197
rect -77 -237 -19 -231
<< nwell >>
rect -263 -369 263 369
<< pmos >>
rect -63 -150 -33 150
rect 33 -150 63 150
<< pdiff >>
rect -125 138 -63 150
rect -125 -138 -113 138
rect -79 -138 -63 138
rect -125 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 125 150
rect 63 -138 79 138
rect 113 -138 125 138
rect 63 -150 125 -138
<< pdiffc >>
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
<< nsubdiff >>
rect -227 299 -131 333
rect 131 299 227 333
rect -227 237 -193 299
rect 193 237 227 299
rect -227 -299 -193 -237
rect 193 -299 227 -237
rect -227 -333 -131 -299
rect 131 -333 227 -299
<< nsubdiffcont >>
rect -131 299 131 333
rect -227 -237 -193 237
rect 193 -237 227 237
rect -131 -333 131 -299
<< poly >>
rect 15 231 81 247
rect 15 197 31 231
rect 65 197 81 231
rect 15 181 81 197
rect -63 150 -33 176
rect 33 150 63 181
rect -63 -181 -33 -150
rect 33 -176 63 -150
rect -81 -197 -15 -181
rect -81 -231 -65 -197
rect -31 -231 -15 -197
rect -81 -247 -15 -231
<< polycont >>
rect 31 197 65 231
rect -65 -231 -31 -197
<< locali >>
rect -227 299 -131 333
rect 131 299 227 333
rect -227 237 -193 299
rect 193 237 227 299
rect 15 197 31 231
rect 65 197 81 231
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
rect -81 -231 -65 -197
rect -31 -231 -15 -197
rect -227 -299 -193 -237
rect 193 -299 227 -237
rect -227 -333 -131 -299
rect 131 -333 227 -299
<< viali >>
rect 31 197 65 231
rect -113 -121 -79 -11
rect -17 11 17 121
rect 79 -121 113 -11
rect -65 -231 -31 -197
<< metal1 >>
rect 19 231 77 237
rect 19 197 31 231
rect 65 197 77 231
rect 19 191 77 197
rect -23 121 23 133
rect -23 11 -17 121
rect 17 11 23 121
rect -119 -11 -73 1
rect -23 -1 23 11
rect -119 -121 -113 -11
rect -79 -121 -73 -11
rect -119 -133 -73 -121
rect 73 -11 119 1
rect 73 -121 79 -11
rect 113 -121 119 -11
rect 73 -133 119 -121
rect -77 -197 -19 -191
rect -77 -231 -65 -197
rect -31 -231 -19 -197
rect -77 -237 -19 -231
<< properties >>
string FIXED_BBOX -210 -316 210 316
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
