** sch_path: /foss/designs/test-xschem/testdp.sch
**.subckt testdp
V8 n GND 0.9
.save i(v8)
Vdd vd GND 1.8
.save i(vdd)
Vc0 c0 GND pulse(1.8 0 0 0 0 5m 10m)
.save i(vc0)
Vc1 c1 GND pulse(1.8 0 0 0 0 10m 20m)
.save i(vc1)
Vc2 c2 GND pulse(1.8 0 0 0 0 20m 40m)
.save i(vc2)
Vc3 c3 GND pulse(1.8 0 0 0 0 40m 80m)
.save i(vc3)
Vc4 c4 GND pulse(1.8 0 0 0 0 80m 160m)
.save i(vc4)
Vc5 c5 GND pulse(1.8 0 0 0 0 160m 320m)
.save i(vc5)
Vc6 c6 GND pulse(1.8 0 0 0 0 320m 640m)
.save i(vc6)
Vc7 c7 GND pulse(1.8 0 0 0 0 640m 1280m)
.save i(vc7)
x1 n GND vd c2 c5 c6 c4 c7 c3 c1 c0 digipot
**** begin user architecture code


.control
save all
*run
tran 1m 1280m 5m
let R = n/i(V8)
plot abs (R)
plot c0 c1+2 c2+4 c3+6 c4+8 c6+10 c7+12
.endc


** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt_mm


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/digipot.sym # of pins=11
** sym_path: /foss/designs/digipot.sym
** sch_path: /foss/designs/digipot.sch
.subckt digipot n gnd vd c2 c5 c6 c4 c7 c3 c1 c0
*.ipin c0
*.ipin c1
*.ipin c2
*.ipin c3
*.ipin c4
*.ipin c5
*.ipin c6
*.ipin c7
*.iopin gnd
*.iopin vd
*.iopin n
XR0 net1 n gnd sky130_fd_pr__res_xhigh_po_0p35 L=22.28 mult=1 m=1
x1 vd c0 gnd net1 gnd tg
XR1 net2 n gnd sky130_fd_pr__res_xhigh_po_0p35 L=10.73 mult=1 m=1
XR2 net3 n gnd sky130_fd_pr__res_xhigh_po_0p35 L=5.48 mult=1 m=1
XR3 net4 n gnd sky130_fd_pr__res_xhigh_po_0p35 L=2.68 mult=1 m=1
XR7 net5 n gnd sky130_fd_pr__res_high_po_0p35 L=0.98 mult=1 m=1
XR6 net6 n gnd sky130_fd_pr__res_high_po_0p35 L=2.07 mult=1 m=1
XR5 net7 n gnd sky130_fd_pr__res_xhigh_po_0p35 L=0.58 mult=1 m=1
XR4 net8 n gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.28 mult=1 m=1
x2 vd c1 gnd net2 gnd tg
x3 vd c2 gnd net3 gnd tg
x4 vd c3 gnd net4 gnd tg
x5 vd c4 gnd net8 gnd tg
x6 vd c5 gnd net7 gnd tg
x7 vd c6 gnd net6 gnd tg
x8 vd c7 gnd net5 gnd tg
.ends


* expanding   symbol:  /foss/designs/tg.sym # of pins=5
** sym_path: /foss/designs/tg.sym
** sch_path: /foss/designs/tg.sch
.subckt tg vd ctrl vgnd A B
*.iopin B
*.iopin A
*.iopin vgnd
*.iopin vd
*.ipin ctrl
x1 vd ctrl nctrl vgnd inverter
XM1 A ctrl B vgnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 A nctrl B vd sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/inverter/xschem_files/inverter.sym # of pins=4
** sym_path: /foss/designs/inverter/xschem_files/inverter.sym
** sch_path: /foss/designs/inverter/xschem_files/inverter.sch
.subckt inverter vd in out gnd
*.ipin in
*.opin out
*.iopin vd
*.iopin gnd
XN0 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XP0 out in vd vd sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
