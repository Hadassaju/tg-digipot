** sch_path: /foss/designs/resistor1.sch
**.subckt resistor1
XR6 net1 net2 net3 sky130_fd_pr__res_high_po_0p35 L=2.07 mult=1 m=1
**.ends
.end
