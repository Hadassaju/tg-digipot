** sch_path: /foss/designs/resistor.sch
**.subckt resistor
XR7 net1 net2 net3 sky130_fd_pr__res_high_po_0p35 L=0.98 mult=1 m=1
**.ends
.end
