magic
tech sky130A
magscale 1 2
timestamp 1698434776
<< pwell >>
rect 460 930 646 1048
rect 752 960 830 1162
<< ndiff >>
rect 852 796 864 908
<< poly >>
rect 1326 658 1432 696
<< metal1 >>
rect 930 1704 1005 1779
rect 930 1364 1005 1664
rect 820 1362 1005 1364
rect 694 1267 1005 1362
rect 694 1257 1004 1267
rect 694 1162 894 1257
rect 1337 1223 1443 1938
rect 1914 1616 1924 1692
rect 2022 1616 2032 1692
rect 1337 1179 1456 1223
rect 381 1056 581 1088
rect 381 918 388 1056
rect 581 930 646 1048
rect 752 960 830 1162
rect 1382 1072 1456 1179
rect 1384 1052 1454 1072
rect 1729 1001 1929 1119
rect 1427 980 1929 1001
rect 756 940 828 960
rect 1260 923 1929 980
rect 1260 920 1480 923
rect 1729 919 1929 923
rect 381 888 581 918
rect 570 744 752 824
rect 830 820 1280 896
rect 1730 792 1930 838
rect 1374 778 1464 780
rect 570 570 650 744
rect 1370 716 1464 778
rect 756 626 826 678
rect 1282 620 1352 678
rect 1000 584 1066 586
rect 1000 570 1200 584
rect 1386 570 1464 716
rect 1564 670 1930 792
rect 1730 638 1930 670
rect 570 490 1466 570
rect 1000 384 1200 490
<< via1 >>
rect 1924 1616 2022 1692
rect 388 918 581 1056
<< metal2 >>
rect 1884 1692 2078 1760
rect 1884 1616 1924 1692
rect 2022 1616 2078 1692
rect 1884 1562 2078 1616
rect 1896 1461 2009 1562
rect 486 1363 2009 1461
rect 486 1115 584 1363
rect 381 1056 584 1115
rect 381 1017 388 1056
rect 385 918 388 1017
rect 581 1017 584 1056
rect 385 908 581 918
rect 385 892 580 908
use sky130_fd_pr__nfet_01v8_A5ES5P  XM1
timestamp 1698428228
transform 1 0 1924 0 1 1757
box 0 0 1 1
use sky130_fd_pr__pfet_01v8_KGAQE3  XM2
timestamp 1698428228
transform 1 0 2293 0 1 3713
box 0 0 1 1
use inverter  inverter_0
timestamp 1698434492
transform -1 0 1294 0 -1 3077
box -793 730 754 1590
use sky130_fd_pr__nfet_01v8_SJYH3Y  sky130_fd_pr__nfet_01v8_SJYH3Y_0
timestamp 1698393312
transform 1 0 791 0 1 808
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_48WM2A  sky130_fd_pr__pfet_01v8_48WM2A_0
timestamp 1698430256
transform 1 0 1370 0 1 863
box -263 -369 263 369
<< labels >>
flabel metal1 1000 384 1200 584 0 FreeSans 256 0 0 0 B
port 4 nsew
flabel metal1 694 1162 894 1362 0 FreeSans 256 0 0 0 ctrl
port 1 nsew
flabel metal1 381 888 581 1088 0 FreeSans 256 0 0 0 vgnd
port 2 nsew
flabel metal1 1730 638 1930 838 0 FreeSans 256 0 0 0 vd
port 0 nsew
flabel metal1 1729 919 1929 1119 0 FreeSans 256 0 0 0 A
port 3 nsew
<< end >>
